-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: Carlos Maytorena
-- 
-- Create Date:    01/06/2020 23:21:32
-- Project Name:   RAM
-- Module Name:    RAM.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity RAM is
   port(D: in STD_LOGIC_VECTOR(8 downto 0);
--		P: inout STD_LOGIC_VECTOR( 15 downto 0);
		Pin: in STD_LOGIC_VECTOR(15 downto 0);
		Pout: out STD_LOGIC_VECTOR(15 downto 0);
		RW,IOM: in STD_LOGIC
		);
end RAM;

architecture arq1 of RAM is

type Ram is array (0 to 511) of STD_LOGIC_VECTOR(15 downto 0);
signal Posicion: Ram:= (x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--30
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--60
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
						x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");

	signal Linea: integer range 0 to 511;

begin

process(D,Pin,Linea)
begin
	Linea<= to_integer(unsigned(D));

	if(IOM = '0') then
		if RW = '1' then
			Posicion(Linea)<= Pin;
		else
			Pout<=Posicion(Linea);
		end if;
	else
		Pout<="ZZZZZZZZZZZZZZZZ";
	end if;

end process;
end arq1;