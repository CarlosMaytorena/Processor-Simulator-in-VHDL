-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: Carlos Maytorena
-- 
-- Create Date:    17/04/2020 11:05:31
-- Project Name:   ROM_Programa
-- Module Name:    ROM_Programa.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity ROM_Programa is
   port(A : in STD_LOGIC_VECTOR(8 downto 0);
		D : out STD_LOGIC_VECTOR(11 downto 0)
		);
end ROM_Programa;

architecture arq1 of ROM_Programa is

	type ROM is array(0 to 511) of STD_LOGIC_VECTOR(11 downto 0);
	constant Programa : ROM :=(x"C10",x"000",x"B04",x"010",x"1D0",x"028",x"BA0",x"010",
							   x"258",x"5D0",x"00F",x"C90",x"010",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",		--30
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",		--60
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
							   x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000");

begin

	D <= Programa(to_integer(unsigned(A)));

end arq1;
