-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: Carlos Maytorena
-- 
-- Create Date:    01/06/2020 20:17:59
-- Project Name:   MemoriadeControl
-- Module Name:    MemoriadeControl.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity MemoriadeControl is
   port(COOP: in STD_LOGIC_VECTOR(11 downto 0);
		Salida: out STD_LOGIC_VECTOR(15 downto 0);
		clk: in STD_LOGIC
		);
end MemoriadeControl;

architecture arq1 of MemoriadeControl is

type Romario is array (0 to 2047) of STD_LOGIC_VECTOR(15 downto 0);

constant Senales: Romario:=(x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--16 SUM mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--21 SUM R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--22 SUM R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--23 SUM R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--25 SUM R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--26 SUM R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--27 SUM R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--29 SUM R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--30 SUM R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--31 SUM R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--32 RES mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--37 RES R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--38 RES R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--39 RES R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--41 RES R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--42 RES R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--43 RES R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--45 RES R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--46 RES R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--47 RES R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--48 MUL mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--50
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",			
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--53 MUL R1,R 
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--54 MUL R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--55 MUL R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--57 MUL R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--58 MUL R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--59 MUL R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--61 MUL R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--62 MUL R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--63 MUL R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--64 DIV mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--69 DIV R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--70 DIV R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--71 DIV R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--73 DIV R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--74 DIV R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--75 DIV R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--77 DIV R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--78 DIV R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--79 DIV R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--80 AND mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--85 AND R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--86 AND R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--87 AND R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--89 AND R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--90 AND R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--91 AND R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--93 AND R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--94 AND R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--95 AND R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--96 OR mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--100
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--101 OR R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--102 OR R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--103 OR R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--105 OR R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--106 OR R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--107 OR R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--109 OR R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--110 OR R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--111 OR R3,#
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0008",x"0000",x"0000",x"0000",x"0000",	--117 NOT R1
							x"4000",x"2800",x"0400",x"0004",x"0000",x"0000",x"0000",x"0000",	--118 NOT R2
							x"4000",x"2800",x"0400",x"0002",x"0000",x"0000",x"0000",x"0000",	--119 NOT R3
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0051",x"0180",	--128 XOR mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",	--133 XOR R1,R
							x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",	--134 XOR R2,R
							x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",	--135 XOR R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0009",x"0000",	--137 XOR R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0005",x"0000",	--138 XOR R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0003",x"0000",	--139 XOR R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0009",x"0000",	--141 XOR R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0005",x"0000",	--142 XOR R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0003",x"0000",	--143 XOR R3,#
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--150
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0041",x"0180",	--160 COMP mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",	--165 COMP R1,R
							x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",	--166 COMP R2,R
							x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",	--167 COMP R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0001",x"0000",	--169 COMP R1,mem 
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0001",x"0000",	--170 COMP R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0001",x"0000",	--171 COMP R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",	
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0001",x"0000",	--173 COMP R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0001",x"0000",	--174 COMP R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0001",x"0000",	--175 COMP R3,#
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0050",x"0180",	--176 MOVE mem,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"0008",x"0000",x"0000",x"0000",x"0000",	--181 MOVE R1,R
							x"4000",x"2800",x"0400",x"0004",x"0000",x"0000",x"0000",x"0000",	--182 MOVE R2,R
							x"4000",x"2800",x"0400",x"0002",x"0000",x"0000",x"0000",x"0000",	--183 MOVE R3,R
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0008",x"0000",	--185 MOVE R1,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0004",x"0000",	--186 MOVE R2,mem
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0010",x"0002",x"0000",	--187 MOVE R3,mem
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0008",x"0000",	--189 MOVE R1,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0004",x"0000",	--190 MOVE R2,#
							x"4000",x"2800",x"0400",x"4000",x"2800",x"0030",x"0002",x"0000",	--191 MOVE R3,#
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0070",x"0008",x"0000",	--193 READ R1,port
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0070",x"0004",x"0000",	--194 READ R2,port
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0070",x"0002",x"0000",	--195 READ R3,port
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--200
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0050",x"0180",x"0000",	--201 WRIT Port,R1
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0050",x"0180",x"0000",	--202 WRIT Port,R2
							x"4000",x"2800",x"0400",x"4000",x"2200",x"0050",x"0180",x"0000",	--203 WRIT Port,R3
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",	--208 JMP dir
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",	--224 JMPL 
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",	--228 JMPE
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",	--232 JMPG 
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",	--240 HALT
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",		--250
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
							x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");

signal PosicionH: STD_LOGIC_VECTOR(10 downto 0);
signal temp_2: STD_LOGIC_VECTOR(2 downto 0);
signal Posicion: integer range 0 to 2047;

begin

process (clk)
	variable temp: unsigned(2 downto 0):= "000";
begin
	if clk'event and clk='1' then	
		temp:= temp+1;	
	end if;
temp_2<= STD_LOGIC_VECTOR(temp);
end process;

PosicionH<=COOP(11 downto 4) & temp_2;
Posicion<= to_integer(unsigned(PosicionH));
Salida <= Senales(Posicion);

end arq1;
